/*
 * Copyright (c) 2024 Andrew Chen
 * SPDX-License-Identifier: Apache-2.0
 */


// Simplified Pong for TinyTapeout
// Testbench to verify behavior
// 640x480 @ 60Hz VGA
// Single paddle + ball

module tb();

endmodule
